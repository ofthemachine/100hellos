module hello_world;

// BEGIN_FRAGLET
initial begin
    $display ("Hello World!");
    $finish;
end
// END_FRAGLET

endmodule